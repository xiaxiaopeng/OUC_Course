---八段数码管显示---
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY DECODER IS
PORT (DATA_IN:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	   DATA_OUT:OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END DECODER;
ARCHITECTURE BHV OF DECODER IS
BEGIN
PROCESS(DATA_IN) 
BEGIN         
		CASE DATA_IN IS 
		    WHEN "0000"=>DATA_OUT<="11000000";
			 WHEN "0001"=>DATA_OUT<="11111001";
			 WHEN "0010"=>DATA_OUT<="10100100"; 
			 WHEN "0011"=>DATA_OUT<="10110000";
			 WHEN "0100"=>DATA_OUT<="10011001";
			 WHEN "0101"=>DATA_OUT<="10010010";
			 WHEN "0110"=>DATA_OUT<="10000010";
			 WHEN "0111"=>DATA_OUT<="11111000";
			 WHEN "1000"=>DATA_OUT<="10000000";
			 WHEN "1001"=>DATA_OUT<="10010000";
			 WHEN OTHERS=>DATA_OUT<="11111111";
			 END CASE;
			 END PROCESS;
END BHV;			 