LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY test5 IS
PORT(				  CLK_50MHz : IN STD_LOGIC;
	CLK_1Hz,CLK_1KHz : OUT STD_LOGIC);
END;
ARCHITECTURE BHV OF test5 IS
SIGNAL Q1 : INTEGER RANGE 0 TO 49999999;
SIGNAL Q2 : INTEGER RANGE 0 TO 199999;
SIGNAL Q3 : INTEGER RANGE 0 TO 9999999;
BEGIN
	PROCESS(CLK_50MHz) BEGIN
		IF CLK_50MHz'EVENT AND CLK_50MHz = '1' THEN
		   -- 1Hz
			IF Q1 < 25000000		THEN CLK_1Hz <= '0'; Q1 <= Q1 + 1;
			ELSIF Q1 < 49999999		THEN CLK_1Hz <= '1'; Q1 <= Q1 + 1;
			ELSE Q1 <= 0;
			END IF;
			-- 1000Hz
			IF Q2 < 25000		THEN CLK_1KHz <= '0'; Q2 <= Q2 + 1;
			ELSIF Q2 < 49999		THEN CLK_1KHz <= '1'; Q2 <= Q2 + 1; 
			ELSE Q2 <= 0;
			END IF;
		END IF;
	END PROCESS;
END;